(* blackbox *)
module SRLC16E (
    output Q,
    Q15,
    input  A0,
    A1,
    A2,
    A3,
    CE,
    CLK,
    D
);
  parameter [15:0] INIT = 16'h0000;
  parameter [0:0] IS_CLK_INVERTED = 1'b0;

  reg [15:0] r = INIT;
  assign Q   = r[{A3, A2, A1, A0}];
  assign Q15 = r[15];
  generate
    begin
      if (IS_CLK_INVERTED) begin
        always @(negedge CLK) if (CE) r <= {r[14:0], D};
      end else begin
        always @(posedge CLK) if (CE) r <= {r[14:0], D};
      end
    end
  endgenerate
endmodule

