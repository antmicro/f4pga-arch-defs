module top (
    output out
);
  assign out = 1;
endmodule  // top
